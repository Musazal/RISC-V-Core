module Control 
	( 
		input [16:0]x, 
		output reg [18:0]y
	);

	always @(*)
	begin
		if (x[6:0] == 'b0110011)
		begin: R_main 
			if (x[16:10] == 'b0000000)
			begin: basic
				case (x[9:7]) 
					0: y = 'b0000000010000000001;
					1: y = 'b0000000010000110001;
					2: y = 'b0000000010000111001;
					3: y = 'b0000000010001101001;
					4: y = 'b0000000010000011001;
					5: y = 'b0000000010000100001;
					6: y = 'b0000000010000010001;
					7: y = 'b0000000010000001001;
					default y = 0;
				endcase
			end
			else if (x[16:10] == 'b0100000)
			begin: sub_sra
				case (x[9:7]) 
					0: y = 'b0000000010001100001;
					5: y = 'b0000000010000101001;
					default: y = 0;
				endcase
			end
			else if (x[16:10] == 'b0000001)
			begin: M_extension
				case (x[9:7]) 
					0: y = 'b0000000010001010001;
					1: y = 'b0000000010001011001;
					2: y = 'b0000000010010100001;
					3: y = 'b0000000010010101001;
					4: y = 'b0000000010001000001;
					5: y = 'b0000000010010110001;
					6: y = 'b0000000010001001001;
					7: y = 'b0000000010010111001;			
					default : y = 0;
				endcase
			end
			else 
				y = 0; 
		end
		else if (x[16:0] == 'b00000010000111011)
			begin: M_W_extension
				y = 'b0000000010010100001;
			end
		else if (x[6:0] == 'b0111011)
		begin: R_word
			if (x[16:10] == 'b0000000)
			begin: basic
				case (x[9:7]) 
					0: y = 'b0000000010001111001;
					1: y = 'b0000000010010001001;
					5: y = 'b0000000010010011001;
					default: y = 0;
				endcase
			end
			else if (x[16:10] == 'b0100000)
			begin: sub_sra 
				case (x[9:7]) 
					0: y = 'b0000000010010000001;
					5: y = 'b0000000010010010001;
					default: y = 0;
				endcase
			end
			else 
				y = 0;
		end
		else if (x[6:0] == 'b0000011)
		begin: Load
			case (x[9:7]) 
				0: y = 'b0000000011000000000;
				1: y = 'b0001000011000000000;
				2: y = 'b0010000011000000000;
				3: y = 'b0011000011000000000;
				4: y = 'b0100000011000000000;
				5: y = 'b0101000011000000000;
				6: y = 'b0110000011000000000;
				default: y = 0;
			endcase
		end
		else if (x[6:0] == 'b0010011)
		begin: I_main
			case (x[9:7]) 
				0: y = 'b0000000011000000001;
				1: begin
					if (x[16:10] == 0) 
						y = 'b0000000011000110001;
					else 
						y = 0;
				end
				2: y = 'b0000000011000111001;
				3: y = 'b0000000011001101001;
				4: y = 'b0000000011000011001;
				5: begin
					if (x[16:10] == 0)
						y = 'b0000000011000100001;
					else 
						y = 'b0000000011000101001;
				end
				6: y = 'b0000000011000010001;
				7: y = 'b0000000011000001001;
				default: y = 0;			
			endcase
		end
		else if (x[6:0] == 'b0011011)
		begin: I_word
			case (x[9:7]) 
				0: y = 'b0000000011001111001;
				1: begin
					if (x[16:10] == 0)
					y = 'b0000000011010001001;
				else
					y = 0;
				end
				5: begin
					if (x[16:10] == 0)
						y = 'b0000000011010010001;
					else 
						y = 'b0000000011010011001;
				end
				default: y = 0;
			endcase
		end
		else if (x[6:0] == 'b1100111)
		begin: jalr
			y = 'b0000100011000000010;
		end
		else if (x[6:0] == 'b0100011)
		begin: Store
			case (x[9:7]) 
				0: y = 'b0000000101000000100;
				1: y = 'b0001000101000000100;
				2: y = 'b0010000101000000100;
				3: y = 'b0011000101000000100;
				default: y = 0;
			endcase
		end
		else if (x[6:0] == 'b1100011)
		begin: Branch
			case (x[9:7]) 
				0: y = 'b1000001000001100000;
				1: y = 'b1000001000001100000;
				4: y = 'b1000001000000111000;
				5: y = 'b1000001000000111000;
				6: y = 'b1000001000001101000;
				7: y = 'b1000001000001101000;
				default: y = 0;
			endcase
		end
		else if (x[6:0] == 'b001011)
		begin:auipc
			y = 'b0000001111100000001;
		end
		else if (x[6:0] == 'b0110111)
		begin:lui
			y = 'b0000001111001110001;
		end
		else if (x[6:0] == 'b1101111)
		begin: jal
			y = 'b0000110011100000010;
		end
		else 
			y = 0;
	end

endmodule 